../../../rtl/rs_monitor.sv