../../../rtl/pre_branch_rtl/data_types.sv