../../../rtl/pre_branch_rtl/broadcast_cdb.sv