../../src/verilog/basic_dmem_model.sv