../../../rtl/instr_fetch_unit.sv