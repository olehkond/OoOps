../../../rtl/instruc_decode.sv