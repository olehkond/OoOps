../../../rtl/pre_branch_rtl/instruc_decode.sv