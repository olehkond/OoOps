../../../src/instructmem.sv