../../../rtl/regfile.sv