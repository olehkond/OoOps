../../../rtl/basic_dmem_model.sv