../../../rtl/OoO_top.sv