../../../rtl/pre_branch_rtl/basic_dmem_model.sv