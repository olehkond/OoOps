../../../rtl/pre_branch_rtl/rs_monitor.sv