../../../rtl/pre_branch_rtl/regfile.sv