../../../rtl/pre_branch_rtl/issue_logic.sv