../../../rtl/load_store_unit.sv