../../../rtl/pre_branch_rtl/alu.sv