../../../rtl/pre_branch_rtl/res_station.sv