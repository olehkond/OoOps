../../../rtl/pre_branch_rtl/OoO_top.sv