../../../rtl/shifter.sv