../../../rtl/branch_unit.sv