../../src/verilog/dmem_read_write_unit.sv