../../../rtl/pre_branch_rtl/dmem_read_write_unit.sv