../../../rtl/branch_pred.sv