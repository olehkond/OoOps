../../../rtl/issue_logic.sv