../../../rtl/fifo.sv