../../../rtl/pre_branch_rtl/fifo.sv