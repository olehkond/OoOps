../../../rtl/broadcast_cdb.sv