../../../rtl/pre_branch_rtl/priority_encoder.sv