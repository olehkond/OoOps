../../../rtl/alu.sv