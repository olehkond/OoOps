../../../rtl/pre_branch_rtl/shifter.sv