../../../rtl/pre_branch_rtl/load_store_unit.sv