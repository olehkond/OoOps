../../../src/datamem.sv