../../../rtl/pre_branch_rtl/alu_br.sv