../../../rtl/res_station.sv