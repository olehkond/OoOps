../../../rtl/priority_encoder.sv