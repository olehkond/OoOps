../../../rtl/data_types.sv