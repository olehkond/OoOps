../../src/verilog/data_types.sv